module PC(
    input [31:0] a,
    output [7:0] b 
);
endmodule