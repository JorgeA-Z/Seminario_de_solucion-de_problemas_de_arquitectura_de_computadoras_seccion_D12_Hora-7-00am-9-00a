module PC(
    input [7:0] a,
    output [7:0] b 
);
endmodule