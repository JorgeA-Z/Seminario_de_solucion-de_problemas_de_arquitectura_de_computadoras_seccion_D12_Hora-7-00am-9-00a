module adder(
    input [7:0] a,
    output [31:0] c);


assign b = 3'b100;

assign c = a + b;
endmodule